CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
21 1Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 18 14 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 537 44 0 3 22
0 8 5 7
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3536 0 0
2
5.89883e-315 5.26354e-315
0
9 2-In AND~
219 365 35 0 3 22
0 3 4 8
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4597 0 0
2
5.89883e-315 5.30499e-315
0
7 Pulser~
4 44 281 0 10 12
0 18 19 2 20 0 0 5 5 4
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3835 0 0
2
5.89883e-315 5.32571e-315
0
2 +V
167 47 10 0 1 3
0 10
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
5.89883e-315 5.34643e-315
0
6 74112~
219 601 184 0 7 32
0 10 7 2 7 10 21 6
0
0 0 4208 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
5616 0 0
2
5.89883e-315 5.3568e-315
0
6 74112~
219 453 189 0 7 32
0 10 8 2 8 10 22 5
0
0 0 4208 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
9323 0 0
2
5.89883e-315 5.36716e-315
0
6 74112~
219 301 187 0 7 32
0 10 3 2 3 10 23 4
0
0 0 4208 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
317 0 0
2
5.89883e-315 5.37752e-315
0
6 74112~
219 145 187 0 7 32
0 10 9 2 9 10 24 3
0
0 0 4208 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3108 0 0
2
5.89883e-315 5.38788e-315
0
9 CC 7-Seg~
183 1019 66 0 18 19
10 17 16 15 14 13 12 11 2 25
0 0 1 1 1 1 1 1 2
0
0 0 21088 0
7 GREENCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4299 0 0
2
5.89883e-315 5.39306e-315
0
6 74LS48
188 846 153 0 14 29
0 6 5 4 3 26 27 11 12 13
14 15 16 17 28
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
5.89883e-315 5.39824e-315
0
36
0 8 2 0 0 4096 0 0 10 19 0 3
566 272
1040 272
1040 102
4 0 3 0 0 12416 0 11 0 0 15 5
814 144
807 144
807 218
195 218
195 151
3 0 4 0 0 12416 0 11 0 0 12 6
814 135
796 135
796 198
337 198
337 107
325 107
2 0 5 0 0 20608 0 11 0 0 8 6
814 126
784 126
784 175
686 175
686 76
477 76
7 1 6 0 0 4224 0 6 11 0 0 4
625 148
773 148
773 117
814 117
4 0 7 0 0 8192 0 6 0 0 7 3
577 166
558 166
558 146
3 2 7 0 0 4224 0 2 6 0 0 3
558 44
558 148
577 148
7 2 5 0 0 0 0 7 2 0 0 3
477 153
477 53
513 53
4 0 8 0 0 4096 0 7 0 0 10 3
429 171
405 171
405 153
2 0 8 0 0 8192 0 7 0 0 11 3
429 153
404 153
404 35
3 1 8 0 0 4224 0 3 2 0 0 2
386 35
513 35
7 2 4 0 0 0 0 8 3 0 0 3
325 151
325 44
341 44
0 1 3 0 0 0 0 0 3 14 0 3
248 151
248 26
341 26
4 0 3 0 0 0 0 8 0 0 15 3
277 169
248 169
248 151
7 2 3 0 0 0 0 9 8 0 0 2
169 151
277 151
4 0 9 0 0 4096 0 9 0 0 21 3
121 169
18 169
18 148
3 0 2 0 0 0 0 7 0 0 19 2
423 162
423 272
3 0 2 0 0 16 0 8 0 0 19 2
271 160
271 272
3 3 2 0 0 4224 0 4 6 0 0 3
68 272
571 272
571 157
3 3 2 0 0 0 0 4 9 0 0 3
68 272
68 160
115 160
1 2 9 0 0 4224 0 1 9 0 0 3
18 26
18 151
121 151
5 0 10 0 0 4096 0 7 0 0 29 2
453 201
453 250
5 0 10 0 0 4096 0 8 0 0 29 2
301 199
301 250
5 0 10 0 0 4096 0 6 0 0 29 2
601 196
601 250
1 0 10 0 0 0 0 6 0 0 29 2
601 121
601 91
1 0 10 0 0 0 0 7 0 0 29 2
453 126
453 91
1 0 10 0 0 0 0 8 0 0 29 2
301 124
301 91
1 0 10 0 0 0 0 9 0 0 29 2
145 124
145 91
1 5 10 0 0 8320 0 5 9 0 0 6
47 19
47 91
674 91
674 250
145 250
145 199
7 7 11 0 0 4224 0 11 10 0 0 3
878 117
1034 117
1034 102
8 6 12 0 0 4224 0 11 10 0 0 3
878 126
1028 126
1028 102
9 5 13 0 0 4224 0 11 10 0 0 3
878 135
1022 135
1022 102
10 4 14 0 0 4224 0 11 10 0 0 3
878 144
1016 144
1016 102
11 3 15 0 0 4224 0 11 10 0 0 3
878 153
1010 153
1010 102
12 2 16 0 0 4224 0 11 10 0 0 3
878 162
1004 162
1004 102
13 1 17 0 0 4224 0 11 10 0 0 3
878 171
998 171
998 102
2
-16 0 0 0 400 0 0 0 0 3 2 1 66
12 Segoe Script
0 0 0 16
156 359 335 400
166 367 324 392
16 GUARIN, AIVAN B.
-16 0 0 0 400 0 0 0 0 3 2 1 2
11 Segoe Print
0 0 0 8
330 357 439 401
340 365 428 393
8 BSCpE-1A
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
